32'h00007033;//  00000000000000000111000000110011;    and r0,r0,r0          h0          
32'h00100093;//  00000000000100000000000010010011;    addi r1,r0, 1         h1 
32'h00200113;//  00000000001000000000000100010011;    addi r2,r0, 2         h2
32'h00308193;//  00000000001100001000000110010011;    addi r3,r1, 3         h4  
32'h00408213;//  00000000010000001000001000010011;    addi r4,r1, 4         h5
32'h00510293;//  00000000010100010000001010010011;    addi r5,r2, 5         h7
32'h00610313;//  00000000011000010000001100010011;    addi r6,r2, 6         h8
32'h00718393;//  00000000011100011000001110010011;    addi r7,r3, 7         hB
32'h00208433;//  00000000001000001000010000110011;    add r8  = r1+r2       h3
32'h404404b3;//  01000000010001000000010010110011;    sub r9  = r8-r4       hfffffffe -2 
32'h00317533;//  00000000001100010111010100110011;    and r10 = r2 & r3     h0
32'h0041e5b3;//  00000000010000011110010110110011;    or  r11 = r3 | r4     h5
32'h02a02823;//  00000010101000000010100000100011;    sw  48(r0)<-- r10     h30 
32'h16802023;//  00010110100000000010000000100011;    sw  352(r0)<-- r8     h160
32'h03002603;//  00000011000000000010011000000011;    lw r12 <-- 48(r0)     for alu result : h30  - for writeback data : h0 
32'h007606B3;//  00000000011101100000011010110011;	  add r13, r12, r7		hB
32'h00311733;//  00000000001100010001011100110011;    sll r14, r2, r3       ALUResult = h20 = r14
32'h408707B3;//  01000000100001110000011110110011;	  sub r15, r14, r8		h1d
32'h00580893;//  00000000010101111000100010010011;	  addi r17, r15, 5  	h22
32'h011909B3;//  00000001000110010000100110110011;	  and r19, r17, r15 	h0